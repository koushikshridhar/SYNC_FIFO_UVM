`include "synchronous_fifo.sv"
`include "top.sv"